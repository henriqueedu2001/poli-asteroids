module digital_circuit (
    
);

endmodule //digital_circuit